library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity PROGRAMA is
    GENERIC( BITS_BUS_DIR   : INTEGER := 8;
             BITS_BUS_DATOS : INTEGER := 15 );
    Port ( BUS_DIR   : in STD_LOGIC_VECTOR  (BITS_BUS_DIR-1 downto 0);
           BUS_DATOS : out STD_LOGIC_VECTOR (BITS_BUS_DATOS-1 downto 0)
           );
end PROGRAMA;

architecture MEMORIA of PROGRAMA is
--CODIGOS DE OPERACION
CONSTANT OP_TR  : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
CONSTANT OP_LI  : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00001";
CONSTANT OP_LWI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00010";
CONSTANT OP_SWI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00011";
CONSTANT OP_ADDI: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00100";
CONSTANT OP_SUBI: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00101";
--SU...
CONSTANT OP_B   : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00110";
CONSTANT OP_CPI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00111";
CONSTANT OP_BEQ : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01000";
CONSTANT OP_BNEQ: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01001";
CONSTANT OP_BLT : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01010";
CONSTANT OP_BLET: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01011";
CONSTANT OP_BGT : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01100";
CONSTANT OP_BGET: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01101";
CONSTANT OP_NOP : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01110";
--CONTINUARA...
--CODIGOS DE FUNCION
CONSTANT FUN_ADD : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
CONSTANT FUN_SUB : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
CONSTANT FUN_AND : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
CONSTANT FUN_OR  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
CONSTANT FUN_XOR : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
CONSTANT FUN_NAND: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
CONSTANT FUN_NOR : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
CONSTANT FUN_XNOR: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";
CONSTANT FUN_CP: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
--CONTINUARA...
CONSTANT SU : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
--REGISTROS
CONSTANT R0 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
CONSTANT R1 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";
CONSTANT R2 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10";
CONSTANT R3 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "11";

TYPE MEM_ROM IS ARRAY( 0 TO 2**BITS_BUS_DIR-1 ) OF STD_LOGIC_VECTOR( BUS_DATOS'RANGE );
CONSTANT MEM_PROG : MEM_ROM := (
    OP_LI&R0&X"01",         --LI R0, #1
    OP_LI&R1&X"07",         --LI R1, #7
    OP_TR&R1&R1&R0&FUN_ADD, --ADD R1, R1, R0
    OP_SWI&R1&X"05",        --SWI R1, 5
    OP_B&SU&X"02",          --B CICLO
    OTHERS => ( OTHERS => '0' )
    --OTHERS => "00000000000000"
    --OTHERS => "000"&X"000"
);

begin

    BUS_DATOS <= MEM_PROG( conv_integer(BUS_DIR) );

end MEMORIA;